`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/18/2025 02:02:41 PM
// Design Name: 
// Module Name: mux2to1
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mux2to1(o, i1, i2, s);
    input [3:0] i1, i2;
    input s;
    output reg [3:0] o;

always @(s or i1 or i2)
begin
    case (s)
        1'b0 : o = i1;
        1'b1 : o = i2;
        default : o = 4'b0;
    endcase
   end
endmodule
